module tb1();
  reg [15:0]i;
  reg [3:0]s; 
  wire out;
  //int a;
  
  mux_16x1 uut(i,s,out);
  
  initial begin
    
    $dumpfile("dump.vcd"); $dumpvars;
    
    i = 16'b0000000000000001; s = 4'b0000; #10;
    i = 16'b0000000000000010; s = 4'b0001; #10;
    i = 16'b0000000000000100; s = 4'b0010; #10;
    i = 16'b0000000000001000; s = 4'b0011; #10;
    i = 16'b0000000000010000; s = 4'b0100; #10;
    i = 16'b0000000000100000; s = 4'b0101; #10;
    i = 16'b0000000001000000; s = 4'b0110; #10;
    i = 16'b0000000010000000; s = 4'b0111; #10;
    i = 16'b0000000100000000; s = 4'b1000; #10;
    i = 16'b0000001000000000; s = 4'b1001; #10;
    i = 16'b0000010000000000; s = 4'b1010; #10;
    i = 16'b0000100000000000; s = 4'b1011; #10;
    i = 16'b0001000000000000; s = 4'b1100; #10;
    i = 16'b0010000000000000; s = 4'b1101; #10;
    i = 16'b0100000000000000; s = 4'b1110; #10;
    i = 16'b1000000000000000; s = 4'b1111; #10;


  end
endmodule